// 1-bit ALU behavioral code
`timescale 1ns/1ps
module alu // Module start declaration
(
  input logic[1:0] a,
  input logic[1:0] b,
  output logic[2:0] c
);
  always@(a or b) 
  begin
    
  end

  
endmodule: alu

